LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY SYSTEM IS
	GENERIC(N: INTEGER := 16);
	PORT(
		DATA 		: INOUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		CLK,RESET,INT	: IN STD_LOGIC
	);
END ENTITY SYSTEM;


ARCHITECTURE SYS_ARCH OF SYSTEM IS


COMPONENT Flag_REG IS
GENERIC (N : INTEGER := 16);
PORT (  IR: IN STD_LOGIC_VECTOR (15 downto 0);
	D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;




COMPONENT REG IS
GENERIC(N : INTEGER := 16);
	PORT(
		CLK,RST	:	IN STD_LOGIC;
		W_EN	:	IN STD_LOGIC;
		D		:	IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		Q		:	OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT DFF IS
	PORT(
		D,CLK,RST	:	IN	STD_LOGIC;
		W_EN		:	IN 	STD_LOGIC;
		Q			:	OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT RAM IS
    GENERIC (
        ADD_WIDTH: INTEGER := 12;
        WRD_WIDTH: INTEGER := 16
    );
    PORT (
        CLK,EN_W,EN_R : IN STD_LOGIC;
	    ADDRESS  : IN STD_LOGIC_VECTOR (ADD_WIDTH-1 DOWNTO 0);
	    DATAIN   : IN STD_LOGIC_VECTOR (WRD_WIDTH-1 DOWNTO 0);
        DATAOUT  : OUT STD_LOGIC_VECTOR (WRD_WIDTH-1 DOWNTO 0)
    );
END COMPONENT;

COMPONENT TRI_STATE_BUFFER IS
    GENERIC(N : INTEGER := 16);
    PORT(
        EN      :   IN  STD_LOGIC;
        INPT    :   IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
        OUTPT   :   OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
    );
END COMPONENT;

COMPONENT ALSU IS
    PORT(
        A,B  : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        S    : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        CIN  : IN STD_LOGIC;
        COUT : OUT STD_LOGIC;
        F    : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        FLAGS  :  OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
    );
END COMPONENT;

COMPONENT M_INS_DEC IS
PORT(IR,FR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	FLAG_OUT: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	CLK,RESET:IN STD_LOGIC;
	OUTPUT: INOUT STD_LOGIC_VECTOR(28 DOWNTO 0));
END COMPONENT;

COMPONENT OP_DECODRS IS
PORT(IR,FR:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	F3:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	IR_BUS_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALU_SELECTORS: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

COMPONENT DECODER_ENABLE IS
	GENERIC (N: INTEGER := 4);
	PORT(
		EN		:	IN STD_LOGIC;
		REG_ADD	:	IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		FOUND	:	OUT STD_LOGIC_VECTOR((2**N)-1 DOWNTO 0)
	);
END COMPONENT;

TYPE GPR IS ARRAY (0 TO 7) OF STD_LOGIC_VECTOR(N-1 DOWNTO 0);
SIGNAL R_data,TI_R : GPR;
SIGNAL TI_SRC,TI_MAR,TI_Y,TI_Z,TI_IR,TI_MDRB,TI_MDRR,TI_MDR : STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL SRC,MAR,Y,Z,IR,MDR : STD_LOGIC_VECTOR (15 DOWNTO 0);
-- SIGNAL SRC_OUT,MAR_OUT,MDR_OUT,Y_OUT,Z_OUT,IR_OUT,MDR_IN : STD_LOGIC_VECTOR (15 DOWNTO 0);
-- SIGNAL SRC_WR,DST_WR,MAR_WR,MDR_WR,Y_WR,Z_WR,IR_WR,SPC_WR: STD_LOGIC;
SIGNAL RAM_IN,RAM_OUT	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL NOT_CLK	:	STD_LOGIC;
SIGNAL MDR_EN	:	STD_LOGIC;
SIGNAL ALU_A,ALU_B,ALU_F	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL ALU_SEL						:	STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL ALU_CIN,ALU_COUT		:	STD_LOGIC;
SIGNAL FLAGIN,FLAGOUT       :   STD_LOGIC_VECTOR (15 DOWNTO 0);
SIGNAL IR_BUS_OUT			:   STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL TRISTATE_ENABLE		: 	STD_LOGIC_VECTOR(28 DOWNTO 0);
SIGNAL CIN_SEL				:	STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL REG_SEL				:	STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL REG_TR_IN_ENABLE,REG_TR_OUT_ENABLE : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL R7_IN_EN,R7_OUT_EN   :	STD_LOGIC;
SIGNAL WRT_DFF,CONTROL_UNIT_RESET	:	STD_LOGIC;
-- SIGNAL TMP_MDR	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
	--GENERAL PURPOSE REGISTERS::
	LP1:FOR i IN 0 TO 6 GENERATE
			TIx: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(REG_TR_IN_ENABLE(i),DATA,TI_R(i));
			Rx: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,REG_TR_IN_ENABLE(i),TI_R(i),R_DATA(i));
			TOx: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(REG_TR_OUT_ENABLE(i),R_DATA(i),DATA);
		END GENERATE;

	TIN_R7: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(R7_IN_EN,DATA,TI_R(7));
	R7: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,R7_IN_EN,TI_R(7),R_DATA(7));
	TOUT_R7: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(R7_OUT_EN,R_DATA(7),DATA);

	TIN_SRC: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(9),DATA,TI_SRC);
	SRC_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(9),TI_SRC,SRC);
	TOUT_SRC: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(26),SRC,DATA);

	TIN_Y: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(0),DATA,TI_Y);
	Y <= TI_Y;	-- JUST FOR THE NAMING CONVENTION
	Y_REG: REG GENERIC MAP (N => 16) PORT MAP(NOT_CLK,RESET,TRISTATE_ENABLE(0),Y,ALU_B);	-- Y outs directly on ALU_B
	-- TOUT_Y: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(RD(9),Y,####ALU####);

	TIN_Z: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(2),ALU_F,TI_Z);	-- ALU_F outs on Z
	Z_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(2),TI_Z,Z);
	TOUT_Z: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(23),Z,DATA);

	TIN_IR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(8),DATA,TI_IR);
	IR_REG: REG GENERIC MAP (N => 16) PORT MAP(NOT_CLK,RESET,TRISTATE_ENABLE(8),TI_IR,IR);			-- REPLACE IR WITH MUHANAD BLACKBOX
	TOUT_IR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(27),IR_BUS_OUT,DATA);

--	TIN_MDRB: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(7),DATA,TI_MDRB);
--	MDRB_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(7),TI_MDRB,TEST1);
--	TOUT_MDRB: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(24),MDR,DATA);

--	TIN_MDRR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(18),RAM_OUT,TEST3);
--	MDRR_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(18),TI_MDRR,TEST2);
--	TOUT_MDRR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(WRT_DFF,MDR,RAM_IN);

	TIN_MDRB: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(7),DATA,TI_MDRB);
	TIN_MDRR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(18),RAM_OUT,TI_MDRR);
	TOUT_MDRB: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(24),MDR,DATA);
	TOUT_MDRR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(WRT_DFF,MDR,RAM_IN);

	TIN_MAR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(TRISTATE_ENABLE(10),DATA,TI_MAR);
	MAR_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(10),TI_MAR,MAR);
--	MAR_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,TRISTATE_ENABLE(10),TI_MAR,MAR);
--	TOUT_MAR: TRI_STATE_BUFFER GENERIC MAP (N => 16) PORT MAP(MAR_EN,MAR,MAR);

--	MAR_EN <= WRT_DFF OR TRISTATE_ENABLE(18);

	WRT_LATCH:	DFF PORT MAP(TRISTATE_ENABLE(19),CLK,RESET,'1',WRT_DFF);


	MDR_EN <= TRISTATE_ENABLE(7) OR TRISTATE_ENABLE(18);

	TI_MDR <= TI_MDRB WHEN TRISTATE_ENABLE(7) ='1'
			ELSE TI_MDRR WHEN TRISTATE_ENABLE(18)='1'
			ELSE (OTHERS => 'Z');


--	MDR <= TEST1 WHEN TRISTATE_ENABLE(7)='1'
--			ELSE TEST2 WHEN TRISTATE_ENABLE(18)='1';

--	TI_MDRR <= RAM_OUT WHEN TRISTATE_ENABLE(18) = '1'
--			ELSE TEST3;

	--REGESTER TO BE SELECTOR BASED ON SRC,DEST
	REG_SEL<= IR(2 DOWNTO 0) WHEN FLAGOUT(5)='1'
 						ELSE	IR(8 DOWNTO 6);

	NOT_CLK <= NOT CLK;
	ALU_A <= DATA;

	R7_IN_EN <= TRISTATE_ENABLE(6) OR REG_TR_IN_ENABLE(7);
	R7_OUT_EN <= TRISTATE_ENABLE(22) OR REG_TR_OUT_ENABLE(7);
	MDR_REG: REG GENERIC MAP (N => 16) PORT MAP(CLK,RESET,MDR_EN,TI_MDR,MDR);


	DECODER_IN_REGISTER: DECODER_ENABLE GENERIC MAP(3) PORT MAP (TRISTATE_ENABLE(3),REG_SEL,REG_TR_IN_ENABLE);
	DECODER_OUT_REGISTER: DECODER_ENABLE GENERIC MAP(3) PORT MAP (TRISTATE_ENABLE(25),REG_SEL,REG_TR_OUT_ENABLE);
	SYS_RAM: RAM GENERIC MAP (WRD_WIDTH => 16,ADD_WIDTH => 12) PORT MAP (NOT_CLK, WRT_DFF, TRISTATE_ENABLE(18), MAR(11 DOWNTO 0), RAM_IN,RAM_OUT);
	--FLAG_REG: REG GENERIC MAP(16) PORT MAP(NOT_CLK,RESET,'1',FLAGIN,FLAGOUT);


	FLAG_REGG: Flag_REG GENERIC MAP(16) PORT MAP(TI_IR,FLAGIN,RESET,CLK,FLAGOUT);


	ALU_OP:	ALSU PORT MAP (ALU_A,ALU_B,ALU_SEL,ALU_CIN,ALU_COUT,ALU_F,FLAGIN(4 DOWNTO 0));
	--OP DECODERS TO HANDLE IR(OFFSET) AND ALU SELECTORS
	ALU_CIN <= CIN_SEL(4);
	ALU_SEL <= CIN_SEL(3 DOWNTO 0);
	OP_ALU_IR: OP_DECODRS PORT MAP(IR,FLAGOUT,TRISTATE_ENABLE(16 DOWNTO 14),IR_BUS_OUT,CIN_SEL);
	CONTROL_UNIT_RESET<=RESET OR INT;
	CONTROL_UNIT: M_INS_DEC PORT MAP (IR,FLAGOUT,FLAGIN(6 DOWNTO 5),CLK,CONTROL_UNIT_RESET,TRISTATE_ENABLE);

END SYS_ARCH;
