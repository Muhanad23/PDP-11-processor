LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY PARTA IS
    PORT(
        A,B : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        S   : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
        CIN : IN STD_LOGIC;
        COUT: OUT STD_LOGIC;
        F   : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END PARTA;

ARCHITECTURE PARTA_FUNC OF PARTA IS
COMPONENT FULL_ADDER IS
    GENERIC (N : INTEGER := 16);
    PORT(
        X,Y  : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
        CIN  : IN STD_LOGIC;
        S    : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
        COUT : OUT STD_LOGIC
    );
END COMPONENT;
    SIGNAL F0,F1,F2,F3,F4,F5,FF,TMPF,NOT_B,B_TCOMP,C_TCOMP: STD_LOGIC_VECTOR (15 DOWNTO 0);
    SIGNAL C0,C1,C2,C3,C4,C5,TMPC,C : STD_LOGIC;
BEGIN
    INC: FULL_ADDER GENERIC MAP (N=>16) PORT MAP(B,"0000000000000000",CIN,F0,C0);        --INCREMENT
    ADC: FULL_ADDER GENERIC MAP (N=>16) PORT MAP(A,B,CIN,F1,C1);                         --ADD WITH CARRY
    SUB: FULL_ADDER GENERIC MAP (N=>16) PORT MAP(A,B_TCOMP,'0',F2,C2);                     --F2=A+(1'S COMPELEMENT OF B)-->(A-B)
    SBC: FULL_ADDER GENERIC MAP (N=>16) PORT MAP(F2,"1111111111111111",'0',F3,C3);        --F3=F2+(1'S COMPELEMENT OF 1)-->(A-B-1)

    --SB: FULL_ADDER GENERIC MAP (N=>16) PORT MAP(TMPF,"0000000000000000",'1',F4,C4);

    u5: FULL_ADDER GENERIC MAP (N=>16) PORT MAP (B,"1111111111111111",'0',F5,C5);        --F5=A+(1'S COMPELEMENT OF 1)-->(A-1)

    u6: FULL_ADDER GENERIC MAP (N=>16) PORT MAP (NOT_B,"0000000000000001",'0',B_TCOMP,C4);        --GET TWO'S COMP
    NOT_B <= NOT B;

		F <= F0 WHEN S="00"
				ELSE F1 WHEN S="01"
				ELSE F3 WHEN S="10" AND CIN='0'
				ELSE F2 WHEN S="10" AND CIN='1'
				ELSE F5 WHEN S="11" AND CIN='0'
				ELSE "0000000000000000";

		COUT <= C0 WHEN S="00"
				ELSE C1 WHEN S="01"
				ELSE C3 WHEN S="10" AND CIN='0'
				ELSE C2 WHEN S="10" AND CIN='1'
				ELSE C5 WHEN S="11" AND CIN='0'
				ELSE '0';

END PARTA_FUNC;
