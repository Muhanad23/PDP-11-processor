LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY CONTROL_UNIT IS
PORT(IR,FR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	FLAG_OUT: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	CLK,RESET:IN STD_LOGIC;
	MICRO_IR:INOUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	M_AR_IN,M_AR_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END ENTITY;

ARCHITECTURE CONT OF CONTROL_UNIT IS
COMPONENT ROM IS
	PORT(
		clk : IN std_logic;
		ADDRESS : IN  std_logic_vector(4 DOWNTO 0);
		DATAOUT : OUT std_logic_vector(17 DOWNTO 0));
END COMPONENT;

COMPONENT DECODING_CIRCUIT IS
PORT(IR,FLAG: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	FLAG_OUT: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	CLK: IN STD_LOGIC;
	NEXT_ADDRESS: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	MICRO_AR: INOUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

COMPONENT TRANSPARENT_REG IS
PORT (D: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

SIGNAL MICRO_AR_IN,MICRO_AR_OUT:STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
	M_AR_OUT<=MICRO_AR_OUT;
	M_AR_IN<=MICRO_AR_IN;
	U0: TRANSPARENT_REG PORT MAP(MICRO_AR_IN,RESET,CLK,MICRO_AR_OUT);
	U1: DECODING_CIRCUIT PORT MAP(IR,FR,FLAG_OUT,CLK,MICRO_IR(17 DOWNTO 13),MICRO_AR_IN);
	U2: ROM PORT MAP(CLK,MICRO_AR_OUT,MICRO_IR);
END ARCHITECTURE;
