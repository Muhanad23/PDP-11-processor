LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY Flag_REG IS
GENERIC (N : INTEGER := 16);
PORT (  IR: IN STD_LOGIC_VECTOR (15 downto 0);
	D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF Flag_REG IS
BEGIN
	PROCESS (CLK)
	BEGIN
		IF (IR(15)='1' and IR(14)='1' and IR(13)='1' and (IR(12))='0') THEN
			Q(5)<='1';
		end if;
		IF (RST='1') THEN
			Q <= (OTHERS => '0');
		ELSIF (RISING_EDGE(CLK)) THEN
			Q <= D;
		END IF;
	end process;
END ARCHITECTURE;	
