LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DFF IS
	PORT(
		D,CLK,RST	:	IN	STD_LOGIC;
		W_EN		:	IN 	STD_LOGIC;
		Q			:	OUT STD_LOGIC
	);
END ENTITY DFF;

ARCHITECTURE DFF_ARCH OF DFF IS
BEGIN
	PROCESS(CLK,RST)
	BEGIN
		IF (RST = '1') THEN
			Q <= '0';
		ELSIF RISING_EDGE(CLK)	THEN
			IF(W_EN = '1')	THEN
			Q <= D;
			END IF;
		END IF;
	END PROCESS;
END DFF_ARCH;