LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY OP_DECODRS IS
PORT(IR,FR:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	F3:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	IR_BUS_OUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	ALU_SELECTORS: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END ENTITY;

ARCHITECTURE OP OF OP_DECODRS IS
SIGNAL BR,ONEOP,F3_SEL:STD_LOGIC;
SIGNAL IR_BUS_OUT_SIG: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL SEL:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL F3_OUT,OP_OUT:STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL OPP: STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
	BR<=IR(15) AND IR(14) AND (NOT IR(13));
	IR_BUS_OUT_SIG<=IR(9)&IR(9)&IR(9)&IR(9)&IR(9)&IR(9)&IR(9 DOWNTO 0);
	ONEOP<=IR(15) AND IR(14) AND IR(13) AND (NOT IR(12));
	F3_SEL<=F3(0) OR F3(1) OR F3(2);

	WITH ONEOP SELECT SEL <=
		IR(15 DOWNTO 12) WHEN '0',
		IR(11 DOWNTO 8) WHEN OTHERS;
	
	WITH BR SELECT IR_BUS_OUT <=
		IR_BUS_OUT_SIG WHEN '1',
		(OTHERS=>'Z') WHEN OTHERS;

	WITH OPP SELECT OP_OUT<=
		--TWO OPERANDS
		"00001" WHEN "00000",
		FR(0)&"0001" WHEN "00001",
		"00010" WHEN "00010" | "00110",
		FR(0)&"0010" WHEN "00011",
		FR(0)&"0110" WHEN "00100",
		FR(0)&"0101" WHEN "00101",
		FR(0)&"0100" WHEN "00111",
		"00000" WHEN "01000",
		--ONE OPERAND
		"10000" WHEN "10000",
		"00011" WHEN "10001",
		"01111" WHEN "10010",
		FR(0)&"0111" WHEN "10011",
		"01000" WHEN "10100",
		"01001" WHEN "10101",
		FR(0)&"1010" WHEN "10110",
		"01011" WHEN "10111",
		"01100" WHEN "11000",
		"01101" WHEN "11001",
		FR(0)&"1110" WHEN "11010",
		(OTHERS=>'Z') WHEN OTHERS;

	OPP(4)<=ONEOP;
	OPP(3 DOWNTO 0)<=SEL;

	WITH F3 SELECT F3_OUT<=
		"10000" WHEN "001",
		"00011" WHEN "010",
		"00001" WHEN "100",
		(OTHERS=>'Z') WHEN OTHERS;

	WITH F3_SEL SELECT ALU_SELECTORS <=
		F3_OUT WHEN '1',
		OP_OUT WHEN OTHERS;
END ARCHITECTURE;