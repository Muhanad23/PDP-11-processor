LIBRARY IEEE;
USE IEEE.std_logic_1164.all;


ENTITY FULL_ADDER IS
    GENERIC (N : INTEGER := 16);
    PORT(
        X,Y  : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
        CIN  : IN STD_LOGIC;
        S    : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
        COUT : OUT STD_LOGIC
    );
END FULL_ADDER;

ARCHITECTURE F_ADDER_FUNC OF FULL_ADDER IS
    COMPONENT HALF_ADDER IS
      PORT(
          X,Y,C : IN STD_LOGIC;
          S,CRY : OUT STD_LOGIC
      );
  END COMPONENT;
SIGNAL CARRY : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
begin
  FX: HALF_ADDER PORT MAP(X(0),Y(0),CIN,S(0),CARRY(0));
  LOOP1: FOR i IN 1 TO N-1 GENERATE
          FI: HALF_ADDER PORT MAP  (X(i),Y(i),CARRY(i-1),S(i),CARRY(i));
    END GENERATE;
    COUT <= CARRY(N-1);
END F_ADDER_FUNC;
