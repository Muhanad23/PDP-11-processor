LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY DECODER IS
GENERIC(N: INTEGER := 3);
PORT (S: IN INTEGER RANGE 0 TO 2**N-1;
	O: OUT STD_LOGIC_VECTOR(2**N-1 DOWNTO 0));
END ENTITY;


ARCHITECTURE BEHAVIOURAL OF DECODER IS
BEGIN
	GEN: FOR I IN 0 To 2**N-1 GENERATE
		O(I) <= '1' WHEN I=S ELSE '0';
	END GENERATE;
END ARCHITECTURE;