LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;

ENTITY DECODER_ENABLE IS
	GENERIC (N: INTEGER := 4);
	PORT(
		EN		:	IN STD_LOGIC;
		REG_ADD	:	IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		FOUND	:	OUT STD_LOGIC_VECTOR((2**N)-1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE DEC_ARCH OF DECODER_ENABLE IS
BEGIN
	GEN: FOR I IN 0 To 2**N-1 GENERATE
		FOUND(I) <= '1' WHEN ((I=to_integer(unsigned(REG_ADD))) AND EN='1')
								ELSE '0';
	END GENERATE;
END ARCHITECTURE;
