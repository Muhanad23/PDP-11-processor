LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE ieee.numeric_std.ALL;

ENTITY M_INS_DEC IS
PORT(IR,FR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	FLAG_OUT: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	CLK,RESET:IN STD_LOGIC;
	OUTPUT: INOUT STD_LOGIC_VECTOR(28 DOWNTO 0));
END ENTITY;

ARCHITECTURE M_INS OF M_INS_DEC IS

COMPONENT CONTROL_UNIT IS
PORT(IR,FR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	FLAG_OUT: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	CLK,RESET:IN STD_LOGIC;
	MICRO_IR:INOUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	M_AR_IN,M_AR_OUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

COMPONENT TRANSPARENT_REG IS
GENERIC (N : INTEGER := 5);
PORT (D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;

COMPONENT DECODER IS
GENERIC(N: INTEGER := 3);
PORT (S: IN INTEGER RANGE 0 TO 2**N-1;
	O: OUT STD_LOGIC_VECTOR(2**N-1 DOWNTO 0));
END COMPONENT;

SIGNAL MIR_IN,MIR_OUT: STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL F1,F2,F3,F4,F5: INTEGER range 0 to 31;
SIGNAL MICRO_AR_IN,MICRO_AR_OUT: STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
	F1<=TO_INTEGER(UNSIGNED(MIR_OUT(12 DOWNTO 10)));
	F2<=TO_INTEGER(UNSIGNED(MIR_OUT(9 DOWNTO 8)));
	F3<=TO_INTEGER(UNSIGNED(MIR_OUT(7 DOWNTO 6)));
	F4<=TO_INTEGER(UNSIGNED(MIR_OUT(5 DOWNTO 3)));
	F5<=TO_INTEGER(UNSIGNED(MIR_OUT(2 DOWNTO 1)));

	U0: CONTROL_UNIT PORT MAP(IR,FR,FLAG_OUT,CLK,RESET,MIR_IN,MICRO_AR_IN,MICRO_AR_OUT);

	U2: TRANSPARENT_REG GENERIC MAP(18)
		PORT MAP(MIR_IN,RESET,CLK,MIR_OUT);

	FF1: DECODER GENERIC MAP(3)
		PORT MAP(F1,OUTPUT(28 DOWNTO 21));
	FF2: DECODER GENERIC MAP(2)
		PORT MAP(F2,OUTPUT(20 DOWNTO 17));
	FF3: DECODER GENERIC MAP(2)
		PORT MAP(F3,OUTPUT(16 DOWNTO 13));
	FF4: DECODER GENERIC MAP(3)
		PORT MAP(F4,OUTPUT(12 DOWNTO 5));
	FF5: DECODER GENERIC MAP(2)
		PORT MAP(F5,OUTPUT(4 DOWNTO 1));
	FF6: OUTPUT(0)<=MIR_OUT(0);

END ARCHITECTURE;
