LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY TRANSPARENT_REG IS
GENERIC (N : INTEGER := 5);
PORT (D: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	RST,CLK: IN STD_LOGIC;
	Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEHAVIOURAL OF TRANSPARENT_REG IS
BEGIN
	PROCESS (CLK)
	BEGIN
		IF (RST='1') THEN
			Q <= (OTHERS => '0');
		ELSIF (RISING_EDGE(CLK)) THEN
			Q <= D;
		END IF;
	END PROCESS;
END ARCHITECTURE;	
